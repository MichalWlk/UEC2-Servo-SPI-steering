`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Michal Walek
// 
// Create Date: 08/02/2024 10:16:12 PM
// Design Name: 
// Module Name: Steering_Y
// Project Name: 
// Target Devices: Basys3
// Tool Versions: 
// Description: Simple divider 100MHz -> 66,67KHz
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Steering_Y(
    input clk,
    input rst,
    input y_val,
    output PWM_y
    );



endmodule