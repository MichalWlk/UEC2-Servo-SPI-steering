//rezultaty musza byc